placerholder
