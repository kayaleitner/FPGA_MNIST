library IEEE;
use IEEE.STD_LOGIC_1164.all;

package denseLayerPkg is

    type array_type is array (natural range<>) of STD_LOGIC_VECTOR;

end denseLayerPkg;

package body denseLayerPkg is 
end denseLayerPkg;