package kernel_pkg is
     type kernel_array_t is array (0 to 8) of integer;
end package kernel_pkg;