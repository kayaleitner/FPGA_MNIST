library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ConvChannel is
end ConvChannel;

architecture beh of ConvChannel is

end beh;
